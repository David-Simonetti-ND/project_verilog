module datapath
(
  input wire [7:0] data ,
  input wire [7:0] key  ,
  input wire clk,
  input wire rst,
  output reg [7:0] encrypted_out
);

    /* something something perform the AES encryption here */

endmodule